//
// VERSAT PROGRAM MEMORY DEFINES
//

