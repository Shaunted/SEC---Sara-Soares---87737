//
// VERSAT REGISTER FILE DEFINES
//

// VERSAT REGISTER FILE ADDRESS WIDTH
`define REGF_ADDR_W 4 //2**4 = 16 registers

// MEMORY MAP
`define R0 `REGF_BASE
`define R1 (`R0+1'b1)
`define R2 (`R1+1'b1)
`define R3 (`R2+1'b1)
`define R4 (`R3+1'b1)
`define R5 (`R4+1'b1)
`define R6 (`R5+1'b1)
`define R7 (`R6+1'b1)
`define R8 (`R7+1'b1)
`define R9 (`R8+1'b1)
`define R10 (`R9+1'b1)
`define R11 (`R10+1'b1)
`define R12 (`R11+1'b1)
`define R13 (`R12+1'b1)
`define R14 (`R13+1'b1)
`define R15 (`R14+1'b1)
